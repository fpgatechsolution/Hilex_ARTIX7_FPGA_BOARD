LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_ARITH.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	LIBRARY xil_defaultlib;
	
	ENTITY hex_seven_seg IS
	PORT(
			osc_clk_in : IN  STD_LOGIC;
						
			KEY_0 :IN STD_LOGIC;
			KEY_1 :IN STD_LOGIC;
			KEY_2 :IN STD_LOGIC;
			KEY_3 :IN STD_LOGIC;
						
			BUZZER:OUT STD_LOGIC;	

			SIG_A : OUT STD_LOGIC;
			SIG_B : OUT STD_LOGIC;
			SIG_C : OUT STD_LOGIC;
			SIG_D : OUT STD_LOGIC;
			SIG_E : OUT STD_LOGIC;
			SIG_F : OUT STD_LOGIC;
			SIG_G : OUT STD_LOGIC;
			SIG_PD: OUT STD_LOGIC;
			SEL_DISP1 : OUT STD_LOGIC;
			SEL_DISP2 : OUT STD_LOGIC;
			SEL_DISP3 : OUT STD_LOGIC;
			SEL_DISP4 : OUT STD_LOGIC;
			
	        LED: OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
			SLIDE_SW: IN  STD_LOGIC_VECTOR (15 DOWNTO 0)
			);
	END hex_seven_seg;
	
	ARCHITECTURE BEHAVIORAL OF hex_seven_seg IS	



SIGNAL RESET:STD_LOGIC;

SIGNAL BCD_VAL_1:STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL BCD_VAL_2:STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL BCD_VAL_3:STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL BCD_VAL_4:STD_LOGIC_VECTOR (3 DOWNTO 0);	

	BEGIN
	
	
	BCD_VAL_1<=SLIDE_SW(3 DOWNTO 0);
	BCD_VAL_2<=SLIDE_SW(7 DOWNTO 4);
	BCD_VAL_3<=SLIDE_SW(11 DOWNTO 8);
	BCD_VAL_4<=SLIDE_SW(15 DOWNTO 12);
	
	LED <=SLIDE_SW;




	RESET <=  KEY_0;
	BUZZER<=  ( KEY_0) OR  ( KEY_1) OR ( KEY_2) OR ( KEY_3);
	
	
	
	
    INST_SEVEN_SEGMENT: ENTITY xil_defaultlib.SEVEN_SEGMENT 
    PORT MAP(
    	CLK_100MHZ =>osc_clk_in ,
    	RESET =>RESET ,
    	SIG_PD =>SIG_PD ,
    	SIG_A =>SIG_A ,
    	SIG_B => SIG_B,
    	SIG_C =>SIG_C ,
    	SIG_D =>SIG_D ,
    	SIG_E =>SIG_E ,
    	SIG_F =>SIG_F ,
    	SIG_G =>SIG_G ,
    	SEL_DISP1 =>SEL_DISP1 ,
    	SEL_DISP2 =>SEL_DISP2 ,
    	SEL_DISP3 =>SEL_DISP3 ,
    	SEL_DISP4 =>SEL_DISP4 ,
    	DATA_DISP_1(3 DOWNTO 0) =>BCD_VAL_1(3 DOWNTO 0) ,
    	DATA_DISP_2(3 DOWNTO 0) =>BCD_VAL_2(3 DOWNTO 0),
    	DATA_DISP_3(3 DOWNTO 0) =>BCD_VAL_3(3 DOWNTO 0) ,
    	DATA_DISP_4(3 DOWNTO 0) =>BCD_VAL_4(3 DOWNTO 0) 
    	);
    
    

	


	END BEHAVIORAL;